library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

entity template is
    Port (
        -- Inputs 
        inv : in std_logic_vector(1 downto 0);
        -- Outputs
        outv : out std_logic_vector(1 downto 0)
    );
end template;

architecture template_arch of template is

begin
    -- Implementation
    
end template_arch;
